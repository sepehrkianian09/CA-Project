module getFour(output [31 : 0] four);
	assign four = 3;
endmodule